module mem_bacnk #(
    parameter ADDR_WIDTH = 16,
    parameter SIZE
) (
    ports
);
    
endmodule